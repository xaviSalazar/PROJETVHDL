LIBRARY       IEEE; 
USE           IEEE.STD_LOGIC_1164.ALL;
use           ieee.std_logic_unsigned.all;
use           IEEE.NUMERIC_STD.all;

entity gestion_anemo is 

port (

--entrees 
clk_50M 			: in std_logic; -- horloge
raz_n           	: in std_logic;	-- reset
in_freq_anemometre  : in std_logic; -- freq du vent
continu				: in std_logic;	-- mode de fonctionnement
start_stop			: in std_logic; -- start/stop
--sorties
data_valid			: out std_logic; -- validation donnee
data_anemometre		: out std_logic_vector (7 downto 0); -- valeur anemo

AffCentaine, AffDizane, AffUnite 		 : out  STD_LOGIC_VECTOR(0 to 6);
clk_1Hz           : out std_logic

);

end gestion_anemo;

architecture behv of gestion_anemo is 
signal valeur_present   : std_logic_vector (25 downto 0):=(others => '0');

signal  debut_periode, fin_periode : std_logic;
signal  periode : std_logic_vector (25 downto 0):=(others => '0');

signal valeur_precedent : std_logic_vector (25 downto 0):=(others => '0');
signal valeur_calcule : std_logic_vector (25 downto 0);

signal centaine, dizaine, unite : std_logic_vector (7 downto 0):=(others => '0');

signal s_data_anemometre		: std_logic_vector (7 downto 0) ;

SIGNAL  count_1Hz      :     unsigned (26 downto 0);

signal s_clk_1Hz           :     std_logic;

BEGIN
-- process pour comptage avec horloge de 50M
process (clk_50M)
begin
	if rising_edge(clk_50M) then
	  if(valeur_present = X"2FAF080") then
	     valeur_present <= (others=>'0');
	  else
	     if(debut_periode = '1') then 
           valeur_present<=valeur_present+X"1";
	    else valeur_present<=valeur_present;
	     end if;
        
	  end if;
	end if;
end process;


div_clk : PROCESS(clk_50M)
begin
if rising_edge(clk_50M) then
if count_1Hz = X"2FAF080" then
centaine <= std_logic_vector(to_unsigned(to_integer( unsigned(s_data_anemometre) / 100), 8));
dizaine  <= std_logic_vector(to_unsigned(to_integer( unsigned (s_data_anemometre) /10  mod 10), 8));
unite    <= std_logic_vector(to_unsigned(to_integer(unsigned (s_data_anemometre) mod 10 ), 8)) ;
s_clk_1Hz<= not s_clk_1Hz;
count_1Hz <= (others => '0');

else
count_1Hz <= count_1Hz + "1";
end IF;
end IF;
end PROCESS div_clk;

clk_1Hz<=s_clk_1Hz;

--deuxieme process
process (in_freq_anemometre)
begin 

	if rising_edge(in_freq_anemometre) then 
        debut_periode <= '1';
		if (valeur_precedent < valeur_present) then
		valeur_calcule <= valeur_present - valeur_precedent;
		elsif (valeur_precedent > valeur_present ) then
        valeur_calcule <= valeur_precedent - valeur_present;
        end if;
        valeur_precedent <= valeur_present;
        
    

     end if;
end process;

s_data_anemometre <=  std_logic_vector(to_unsigned( to_integer( 50000000 / unsigned (valeur_calcule)) ,8 ) );
data_anemometre <= s_data_anemometre;

--centaine <= std_logic_vector(to_unsigned(to_integer( unsigned(s_data_anemometre) / 100), 8));
--dizaine  <= std_logic_vector(to_unsigned(to_integer( unsigned (s_data_anemometre) /10  mod 10), 8));
--unite    <= std_logic_vector(to_unsigned(to_integer(unsigned (s_data_anemometre) mod 10 ), 8)) ;


AffCentaine <=  "0000001" when centaine =X"00"   else
                "1001111" when centaine =X"01"   else
                "0010010" when centaine =X"02"   else
                "0000110" when centaine =X"03"   else
                "1001100" when centaine =X"04"   else
                "0100100" when centaine =X"05"   else
                "0100000" when centaine =X"06"   else
                "0001111" when centaine =X"07"   else
                "0000000" when centaine =X"08"   else
                "0000100" when centaine =X"09"   else
                "1111111";
                
AffDizane <=    "0000001" when dizaine =X"00"   else
                "1001111" when dizaine =X"01"   else
                "0010010" when dizaine =X"02"   else
                "0000110" when dizaine =X"03"   else
                "1001100" when dizaine =X"04"   else
                "0100100" when dizaine =X"05"   else
                "0100000" when dizaine =X"06"   else
                "0001111" when dizaine =X"07"   else
                "0000000" when dizaine =X"08"   else
                "0000100" when dizaine =X"09"   else
                "1111111";
                
AffUnite <=     "0000001" when unite =X"00"   else
                "1001111" when unite =X"01"   else
                "0010010" when unite =X"02"   else
                "0000110" when unite =X"03"   else
                "1001100" when unite =X"04"   else
                "0100100" when unite =X"05"   else
                "0100000" when unite =X"06"   else
                "0001111" when unite =X"07"   else
                "0000000" when unite =X"08"   else
                "0000100" when unite =X"09"   else
                "1111111";             

END behv;








--LIBRARY       IEEE; 
--USE           IEEE.STD_LOGIC_1164.ALL;
--use           ieee.std_logic_unsigned.all;
--use           IEEE.NUMERIC_STD.all;
--
--entity gestion_anemo is 
--
--port (
--
----entrees 
--clk_50M 			: in std_logic; -- horloge
--raz_n           	: in std_logic;	-- reset
--in_freq_anemometre  : in std_logic; -- freq du vent
--continu				: in std_logic;	-- mode de fonctionnement
--start_stop			: in std_logic; -- start/stop
----sorties
--data_valid			: out std_logic; -- validation donnee
--data_anemometre		: out std_logic_vector (7 downto 0); -- valeur anemo
--
--AffCentaine, AffDizane, AffUnite 		 : out  STD_LOGIC_VECTOR(0 to 6);
--clk_200Hz           : out std_logic
--
--);
--
--end gestion_anemo;
--
--architecture behv of gestion_anemo is 
--signal valeur_present   : std_logic_vector (25 downto 0):=(others => '0');
--
--signal  etatHaut : std_logic_vector (25 downto 0):=(others => '0');
--signal  etatBas : std_logic_vector (25 downto 0):=(others => '0');
--signal  etat : std_logic;
--signal periode : std_logic_vector (25 downto 0):=(others => '0');
--
----signal  etatHaut : std_logic;
----signal  etatBas : std_logic;
----signal  variable1 : std_logic_vector (25 downto 0):=(others => '0');
----signal  variable2 : std_logic_vector (25 downto 0):=(others => '0');
----signal  period2 : std_logic_vector (25 downto 0):=(others => '0');
----signal  period1 : std_logic_vector (25 downto 0):=(others => '0');
--
--
--signal valeur_precedent : std_logic_vector (25 downto 0):=(others => '0');
--signal valeur_calcule : std_logic_vector (25 downto 0);
--
--signal centaine, dizaine, unite : std_logic_vector (7 downto 0):=(others => '0');
--
--signal s_data_anemometre		: std_logic_vector (7 downto 0) ;
--
--SIGNAL  count_200Hz      :     unsigned (26 downto 0);
--signal s_clk_200Hz           :     std_logic;
--
--BEGIN
---- process pour comptage avec horloge de 50M
--process (clk_50M)
--begin
--	if rising_edge(clk_50M) then
----	-------------------------------------------------------
----				if(etatHaut = '1' and etatBas = '0') then  
----					variable1 <= variable1+x"1";
----				end if;
----				
----				if(etatHaut = '0' and etatBas = '1') then  
----					variable2 <= variable2+x"1";
----				end if;
----		
----	---------------------------------------------------------
--	    if(etatHaut = X"2FAF080") then etatHaut <= (others => '0');
--	    else
--	       if(etatBas = X"2FAF080") then etatBas <= (others => '0');
--           end if;
--        end if;
--
--	    if(etat='0') then etatBas <= etatBas + X"1";
--	    else
--	       if(etat='1') then etatHaut <= etatHaut + X"1";
--		--valeur_present <= valeur_present + X"1";
--	       end if;
--	     end if;
--
--        if count_200Hz = X"7A120" then
--         s_clk_200Hz<= not s_clk_200Hz;
--         count_200Hz <= (others => '0');
--        else
--          count_200Hz <= count_200Hz + "1";
--        end if; 
---------------------------------------------------------------------
--	end if;
--end process;
--
--clk_200Hz<=s_clk_200Hz;
--
----deuxieme process
--process (in_freq_anemometre)
--begin 
---------------------------------------------------------------
----if rising_edge(in_freq_anemometre) then
----variable1 <= (others=>'0');
----period2 <= variable2;
----etatHaut <= '1';
----etatBas <= '0';
----
----else 
----if falling_edge(in_freq_anemometre) then
------
----variable2 <= (others=>'0');
----period1 <= variable1;
----etatHaut <= '0';
----etatBas <= '1';
----end if;
----end if;
------------------------------------------------------------------
--	if rising_edge(in_freq_anemometre) then
--        etat<='1';
--    else
--        if falling_edge(in_freq_anemometre) then
--        etat<='0';
--        else etat<='X';
--        end if;
--     end if;
--	--	if (valeur_precedent < valeur_present) then
--	--	valeur_calcule <= valeur_present - valeur_precedent;
--	--	elsif (valeur_precedent > valeur_present ) then
--    --    valeur_calcule <= valeur_precedent - valeur_present;
--    --    end if;
--    --    valeur_precedent <= valeur_present;
--    -- end if;
--    if(etatHaut /= X"0" and etatBas /= X"0") then 
--    valeur_calcule <= etatBas + etatHaut;
--     etatHaut <= (others => '0');
--    etatBas <= (others => '0');  
--    end if;  
--end process;
--
--s_data_anemometre <=  std_logic_vector(to_unsigned( to_integer( 50000000 / unsigned (valeur_calcule)) ,8 ) );
--data_anemometre <= s_data_anemometre;
--
--centaine <= std_logic_vector(to_unsigned(to_integer( unsigned(s_data_anemometre) / 100), 8));
--dizaine  <= std_logic_vector(to_unsigned(to_integer( unsigned (s_data_anemometre) /10  mod 10), 8));
--unite    <= std_logic_vector(to_unsigned(to_integer(unsigned (s_data_anemometre) mod 10 ), 8)) ;
--
--AffCentaine <=  "0000001" when centaine =X"00"   else
--                "1001111" when centaine =X"01"   else
--                "0010010" when centaine =X"02"   else
--                "0000110" when centaine =X"03"   else
--                "1001100" when centaine =X"04"   else
--                "0100100" when centaine =X"05"   else
--                "0100000" when centaine =X"06"   else
--                "0001111" when centaine =X"07"   else
--                "0000000" when centaine =X"08"   else
--                "0000100" when centaine =X"09"   else
--                "1111111";
--                
--AffDizane <=    "0000001" when dizaine =X"00"   else
--                "1001111" when dizaine =X"01"   else
--                "0010010" when dizaine =X"02"   else
--                "0000110" when dizaine =X"03"   else
--                "1001100" when dizaine =X"04"   else
--                "0100100" when dizaine =X"05"   else
--                "0100000" when dizaine =X"06"   else
--                "0001111" when dizaine =X"07"   else
--                "0000000" when dizaine =X"08"   else
--                "0000100" when dizaine =X"09"   else
--                "1111111";
--                
--AffUnite <=     "0000001" when unite =X"00"   else
--                "1001111" when unite =X"01"   else
--                "0010010" when unite =X"02"   else
--                "0000110" when unite =X"03"   else
--                "1001100" when unite =X"04"   else
--                "0100100" when unite =X"05"   else
--                "0100000" when unite =X"06"   else
--                "0001111" when unite =X"07"   else
--                "0000000" when unite =X"08"   else
--                "0000100" when unite =X"09"   else
--                "1111111";
--               
--
--END behv;


